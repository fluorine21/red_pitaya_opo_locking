//Sine wave lookup table with 1024 points
//Regenerate using sine_wave_rom_gen.m

import opo_package::*;

module sine_lut(
 input wire [sine_lut_width-1:0] addr,
output reg [word_width-1:0] data
);

always @ * begin

case(addr)

10'h0000 : data = 16'h0000;
10'h0001 : data = 16'h00C9;
10'h0002 : data = 16'h0192;
10'h0003 : data = 16'h025B;
10'h0004 : data = 16'h0324;
10'h0005 : data = 16'h03ED;
10'h0006 : data = 16'h04B6;
10'h0007 : data = 16'h057F;
10'h0008 : data = 16'h0648;
10'h0009 : data = 16'h0711;
10'h000A : data = 16'h07D9;
10'h000B : data = 16'h08A2;
10'h000C : data = 16'h096A;
10'h000D : data = 16'h0A33;
10'h000E : data = 16'h0AFB;
10'h000F : data = 16'h0BC4;
10'h0010 : data = 16'h0C8C;
10'h0011 : data = 16'h0D54;
10'h0012 : data = 16'h0E1C;
10'h0013 : data = 16'h0EE3;
10'h0014 : data = 16'h0FAB;
10'h0015 : data = 16'h1072;
10'h0016 : data = 16'h113A;
10'h0017 : data = 16'h1201;
10'h0018 : data = 16'h12C8;
10'h0019 : data = 16'h138F;
10'h001A : data = 16'h1455;
10'h001B : data = 16'h151C;
10'h001C : data = 16'h15E2;
10'h001D : data = 16'h16A8;
10'h001E : data = 16'h176E;
10'h001F : data = 16'h1833;
10'h0020 : data = 16'h18F9;
10'h0021 : data = 16'h19BE;
10'h0022 : data = 16'h1A82;
10'h0023 : data = 16'h1B47;
10'h0024 : data = 16'h1C0B;
10'h0025 : data = 16'h1CCF;
10'h0026 : data = 16'h1D93;
10'h0027 : data = 16'h1E57;
10'h0028 : data = 16'h1F1A;
10'h0029 : data = 16'h1FDD;
10'h002A : data = 16'h209F;
10'h002B : data = 16'h2161;
10'h002C : data = 16'h2223;
10'h002D : data = 16'h22E5;
10'h002E : data = 16'h23A6;
10'h002F : data = 16'h2467;
10'h0030 : data = 16'h2528;
10'h0031 : data = 16'h25E8;
10'h0032 : data = 16'h26A8;
10'h0033 : data = 16'h2767;
10'h0034 : data = 16'h2826;
10'h0035 : data = 16'h28E5;
10'h0036 : data = 16'h29A3;
10'h0037 : data = 16'h2A61;
10'h0038 : data = 16'h2B1F;
10'h0039 : data = 16'h2BDC;
10'h003A : data = 16'h2C99;
10'h003B : data = 16'h2D55;
10'h003C : data = 16'h2E11;
10'h003D : data = 16'h2ECC;
10'h003E : data = 16'h2F87;
10'h003F : data = 16'h3041;
10'h0040 : data = 16'h30FB;
10'h0041 : data = 16'h31B5;
10'h0042 : data = 16'h326E;
10'h0043 : data = 16'h3326;
10'h0044 : data = 16'h33DF;
10'h0045 : data = 16'h3496;
10'h0046 : data = 16'h354D;
10'h0047 : data = 16'h3604;
10'h0048 : data = 16'h36BA;
10'h0049 : data = 16'h376F;
10'h004A : data = 16'h3824;
10'h004B : data = 16'h38D9;
10'h004C : data = 16'h398C;
10'h004D : data = 16'h3A40;
10'h004E : data = 16'h3AF2;
10'h004F : data = 16'h3BA5;
10'h0050 : data = 16'h3C56;
10'h0051 : data = 16'h3D07;
10'h0052 : data = 16'h3DB8;
10'h0053 : data = 16'h3E68;
10'h0054 : data = 16'h3F17;
10'h0055 : data = 16'h3FC5;
10'h0056 : data = 16'h4073;
10'h0057 : data = 16'h4121;
10'h0058 : data = 16'h41CE;
10'h0059 : data = 16'h427A;
10'h005A : data = 16'h4325;
10'h005B : data = 16'h43D0;
10'h005C : data = 16'h447A;
10'h005D : data = 16'h4524;
10'h005E : data = 16'h45CD;
10'h005F : data = 16'h4675;
10'h0060 : data = 16'h471C;
10'h0061 : data = 16'h47C3;
10'h0062 : data = 16'h4869;
10'h0063 : data = 16'h490F;
10'h0064 : data = 16'h49B4;
10'h0065 : data = 16'h4A58;
10'h0066 : data = 16'h4AFB;
10'h0067 : data = 16'h4B9D;
10'h0068 : data = 16'h4C3F;
10'h0069 : data = 16'h4CE0;
10'h006A : data = 16'h4D81;
10'h006B : data = 16'h4E20;
10'h006C : data = 16'h4EBF;
10'h006D : data = 16'h4F5D;
10'h006E : data = 16'h4FFB;
10'h006F : data = 16'h5097;
10'h0070 : data = 16'h5133;
10'h0071 : data = 16'h51CE;
10'h0072 : data = 16'h5268;
10'h0073 : data = 16'h5302;
10'h0074 : data = 16'h539B;
10'h0075 : data = 16'h5432;
10'h0076 : data = 16'h54C9;
10'h0077 : data = 16'h5560;
10'h0078 : data = 16'h55F5;
10'h0079 : data = 16'h568A;
10'h007A : data = 16'h571D;
10'h007B : data = 16'h57B0;
10'h007C : data = 16'h5842;
10'h007D : data = 16'h58D3;
10'h007E : data = 16'h5964;
10'h007F : data = 16'h59F3;
10'h0080 : data = 16'h5A82;
10'h0081 : data = 16'h5B0F;
10'h0082 : data = 16'h5B9C;
10'h0083 : data = 16'h5C28;
10'h0084 : data = 16'h5CB3;
10'h0085 : data = 16'h5D3E;
10'h0086 : data = 16'h5DC7;
10'h0087 : data = 16'h5E4F;
10'h0088 : data = 16'h5ED7;
10'h0089 : data = 16'h5F5D;
10'h008A : data = 16'h5FE3;
10'h008B : data = 16'h6068;
10'h008C : data = 16'h60EB;
10'h008D : data = 16'h616E;
10'h008E : data = 16'h61F0;
10'h008F : data = 16'h6271;
10'h0090 : data = 16'h62F1;
10'h0091 : data = 16'h6370;
10'h0092 : data = 16'h63EE;
10'h0093 : data = 16'h646C;
10'h0094 : data = 16'h64E8;
10'h0095 : data = 16'h6563;
10'h0096 : data = 16'h65DD;
10'h0097 : data = 16'h6656;
10'h0098 : data = 16'h66CF;
10'h0099 : data = 16'h6746;
10'h009A : data = 16'h67BC;
10'h009B : data = 16'h6832;
10'h009C : data = 16'h68A6;
10'h009D : data = 16'h6919;
10'h009E : data = 16'h698B;
10'h009F : data = 16'h69FD;
10'h00A0 : data = 16'h6A6D;
10'h00A1 : data = 16'h6ADC;
10'h00A2 : data = 16'h6B4A;
10'h00A3 : data = 16'h6BB7;
10'h00A4 : data = 16'h6C23;
10'h00A5 : data = 16'h6C8E;
10'h00A6 : data = 16'h6CF8;
10'h00A7 : data = 16'h6D61;
10'h00A8 : data = 16'h6DC9;
10'h00A9 : data = 16'h6E30;
10'h00AA : data = 16'h6E96;
10'h00AB : data = 16'h6EFB;
10'h00AC : data = 16'h6F5E;
10'h00AD : data = 16'h6FC1;
10'h00AE : data = 16'h7022;
10'h00AF : data = 16'h7083;
10'h00B0 : data = 16'h70E2;
10'h00B1 : data = 16'h7140;
10'h00B2 : data = 16'h719D;
10'h00B3 : data = 16'h71F9;
10'h00B4 : data = 16'h7254;
10'h00B5 : data = 16'h72AE;
10'h00B6 : data = 16'h7307;
10'h00B7 : data = 16'h735E;
10'h00B8 : data = 16'h73B5;
10'h00B9 : data = 16'h740A;
10'h00BA : data = 16'h745F;
10'h00BB : data = 16'h74B2;
10'h00BC : data = 16'h7504;
10'h00BD : data = 16'h7555;
10'h00BE : data = 16'h75A5;
10'h00BF : data = 16'h75F3;
10'h00C0 : data = 16'h7641;
10'h00C1 : data = 16'h768D;
10'h00C2 : data = 16'h76D8;
10'h00C3 : data = 16'h7722;
10'h00C4 : data = 16'h776B;
10'h00C5 : data = 16'h77B3;
10'h00C6 : data = 16'h77FA;
10'h00C7 : data = 16'h783F;
10'h00C8 : data = 16'h7884;
10'h00C9 : data = 16'h78C7;
10'h00CA : data = 16'h7909;
10'h00CB : data = 16'h794A;
10'h00CC : data = 16'h7989;
10'h00CD : data = 16'h79C8;
10'h00CE : data = 16'h7A05;
10'h00CF : data = 16'h7A41;
10'h00D0 : data = 16'h7A7C;
10'h00D1 : data = 16'h7AB6;
10'h00D2 : data = 16'h7AEE;
10'h00D3 : data = 16'h7B26;
10'h00D4 : data = 16'h7B5C;
10'h00D5 : data = 16'h7B91;
10'h00D6 : data = 16'h7BC5;
10'h00D7 : data = 16'h7BF8;
10'h00D8 : data = 16'h7C29;
10'h00D9 : data = 16'h7C59;
10'h00DA : data = 16'h7C88;
10'h00DB : data = 16'h7CB6;
10'h00DC : data = 16'h7CE3;
10'h00DD : data = 16'h7D0E;
10'h00DE : data = 16'h7D39;
10'h00DF : data = 16'h7D62;
10'h00E0 : data = 16'h7D89;
10'h00E1 : data = 16'h7DB0;
10'h00E2 : data = 16'h7DD5;
10'h00E3 : data = 16'h7DFA;
10'h00E4 : data = 16'h7E1D;
10'h00E5 : data = 16'h7E3E;
10'h00E6 : data = 16'h7E5F;
10'h00E7 : data = 16'h7E7E;
10'h00E8 : data = 16'h7E9C;
10'h00E9 : data = 16'h7EB9;
10'h00EA : data = 16'h7ED5;
10'h00EB : data = 16'h7EEF;
10'h00EC : data = 16'h7F09;
10'h00ED : data = 16'h7F21;
10'h00EE : data = 16'h7F37;
10'h00EF : data = 16'h7F4D;
10'h00F0 : data = 16'h7F61;
10'h00F1 : data = 16'h7F74;
10'h00F2 : data = 16'h7F86;
10'h00F3 : data = 16'h7F97;
10'h00F4 : data = 16'h7FA6;
10'h00F5 : data = 16'h7FB4;
10'h00F6 : data = 16'h7FC1;
10'h00F7 : data = 16'h7FCD;
10'h00F8 : data = 16'h7FD8;
10'h00F9 : data = 16'h7FE1;
10'h00FA : data = 16'h7FE9;
10'h00FB : data = 16'h7FF0;
10'h00FC : data = 16'h7FF5;
10'h00FD : data = 16'h7FF9;
10'h00FE : data = 16'h7FFD;
10'h00FF : data = 16'h7FFE;
10'h0100 : data = 16'h7FFF;
10'h0101 : data = 16'h7FFE;
10'h0102 : data = 16'h7FFD;
10'h0103 : data = 16'h7FF9;
10'h0104 : data = 16'h7FF5;
10'h0105 : data = 16'h7FF0;
10'h0106 : data = 16'h7FE9;
10'h0107 : data = 16'h7FE1;
10'h0108 : data = 16'h7FD8;
10'h0109 : data = 16'h7FCD;
10'h010A : data = 16'h7FC1;
10'h010B : data = 16'h7FB4;
10'h010C : data = 16'h7FA6;
10'h010D : data = 16'h7F97;
10'h010E : data = 16'h7F86;
10'h010F : data = 16'h7F74;
10'h0110 : data = 16'h7F61;
10'h0111 : data = 16'h7F4D;
10'h0112 : data = 16'h7F37;
10'h0113 : data = 16'h7F21;
10'h0114 : data = 16'h7F09;
10'h0115 : data = 16'h7EEF;
10'h0116 : data = 16'h7ED5;
10'h0117 : data = 16'h7EB9;
10'h0118 : data = 16'h7E9C;
10'h0119 : data = 16'h7E7E;
10'h011A : data = 16'h7E5F;
10'h011B : data = 16'h7E3E;
10'h011C : data = 16'h7E1D;
10'h011D : data = 16'h7DFA;
10'h011E : data = 16'h7DD5;
10'h011F : data = 16'h7DB0;
10'h0120 : data = 16'h7D89;
10'h0121 : data = 16'h7D62;
10'h0122 : data = 16'h7D39;
10'h0123 : data = 16'h7D0E;
10'h0124 : data = 16'h7CE3;
10'h0125 : data = 16'h7CB6;
10'h0126 : data = 16'h7C88;
10'h0127 : data = 16'h7C59;
10'h0128 : data = 16'h7C29;
10'h0129 : data = 16'h7BF8;
10'h012A : data = 16'h7BC5;
10'h012B : data = 16'h7B91;
10'h012C : data = 16'h7B5C;
10'h012D : data = 16'h7B26;
10'h012E : data = 16'h7AEE;
10'h012F : data = 16'h7AB6;
10'h0130 : data = 16'h7A7C;
10'h0131 : data = 16'h7A41;
10'h0132 : data = 16'h7A05;
10'h0133 : data = 16'h79C8;
10'h0134 : data = 16'h7989;
10'h0135 : data = 16'h794A;
10'h0136 : data = 16'h7909;
10'h0137 : data = 16'h78C7;
10'h0138 : data = 16'h7884;
10'h0139 : data = 16'h783F;
10'h013A : data = 16'h77FA;
10'h013B : data = 16'h77B3;
10'h013C : data = 16'h776B;
10'h013D : data = 16'h7722;
10'h013E : data = 16'h76D8;
10'h013F : data = 16'h768D;
10'h0140 : data = 16'h7641;
10'h0141 : data = 16'h75F3;
10'h0142 : data = 16'h75A5;
10'h0143 : data = 16'h7555;
10'h0144 : data = 16'h7504;
10'h0145 : data = 16'h74B2;
10'h0146 : data = 16'h745F;
10'h0147 : data = 16'h740A;
10'h0148 : data = 16'h73B5;
10'h0149 : data = 16'h735E;
10'h014A : data = 16'h7307;
10'h014B : data = 16'h72AE;
10'h014C : data = 16'h7254;
10'h014D : data = 16'h71F9;
10'h014E : data = 16'h719D;
10'h014F : data = 16'h7140;
10'h0150 : data = 16'h70E2;
10'h0151 : data = 16'h7083;
10'h0152 : data = 16'h7022;
10'h0153 : data = 16'h6FC1;
10'h0154 : data = 16'h6F5E;
10'h0155 : data = 16'h6EFB;
10'h0156 : data = 16'h6E96;
10'h0157 : data = 16'h6E30;
10'h0158 : data = 16'h6DC9;
10'h0159 : data = 16'h6D61;
10'h015A : data = 16'h6CF8;
10'h015B : data = 16'h6C8E;
10'h015C : data = 16'h6C23;
10'h015D : data = 16'h6BB7;
10'h015E : data = 16'h6B4A;
10'h015F : data = 16'h6ADC;
10'h0160 : data = 16'h6A6D;
10'h0161 : data = 16'h69FD;
10'h0162 : data = 16'h698B;
10'h0163 : data = 16'h6919;
10'h0164 : data = 16'h68A6;
10'h0165 : data = 16'h6832;
10'h0166 : data = 16'h67BC;
10'h0167 : data = 16'h6746;
10'h0168 : data = 16'h66CF;
10'h0169 : data = 16'h6656;
10'h016A : data = 16'h65DD;
10'h016B : data = 16'h6563;
10'h016C : data = 16'h64E8;
10'h016D : data = 16'h646C;
10'h016E : data = 16'h63EE;
10'h016F : data = 16'h6370;
10'h0170 : data = 16'h62F1;
10'h0171 : data = 16'h6271;
10'h0172 : data = 16'h61F0;
10'h0173 : data = 16'h616E;
10'h0174 : data = 16'h60EB;
10'h0175 : data = 16'h6068;
10'h0176 : data = 16'h5FE3;
10'h0177 : data = 16'h5F5D;
10'h0178 : data = 16'h5ED7;
10'h0179 : data = 16'h5E4F;
10'h017A : data = 16'h5DC7;
10'h017B : data = 16'h5D3E;
10'h017C : data = 16'h5CB3;
10'h017D : data = 16'h5C28;
10'h017E : data = 16'h5B9C;
10'h017F : data = 16'h5B0F;
10'h0180 : data = 16'h5A82;
10'h0181 : data = 16'h59F3;
10'h0182 : data = 16'h5964;
10'h0183 : data = 16'h58D3;
10'h0184 : data = 16'h5842;
10'h0185 : data = 16'h57B0;
10'h0186 : data = 16'h571D;
10'h0187 : data = 16'h568A;
10'h0188 : data = 16'h55F5;
10'h0189 : data = 16'h5560;
10'h018A : data = 16'h54C9;
10'h018B : data = 16'h5432;
10'h018C : data = 16'h539B;
10'h018D : data = 16'h5302;
10'h018E : data = 16'h5268;
10'h018F : data = 16'h51CE;
10'h0190 : data = 16'h5133;
10'h0191 : data = 16'h5097;
10'h0192 : data = 16'h4FFB;
10'h0193 : data = 16'h4F5D;
10'h0194 : data = 16'h4EBF;
10'h0195 : data = 16'h4E20;
10'h0196 : data = 16'h4D81;
10'h0197 : data = 16'h4CE0;
10'h0198 : data = 16'h4C3F;
10'h0199 : data = 16'h4B9D;
10'h019A : data = 16'h4AFB;
10'h019B : data = 16'h4A58;
10'h019C : data = 16'h49B4;
10'h019D : data = 16'h490F;
10'h019E : data = 16'h4869;
10'h019F : data = 16'h47C3;
10'h01A0 : data = 16'h471C;
10'h01A1 : data = 16'h4675;
10'h01A2 : data = 16'h45CD;
10'h01A3 : data = 16'h4524;
10'h01A4 : data = 16'h447A;
10'h01A5 : data = 16'h43D0;
10'h01A6 : data = 16'h4325;
10'h01A7 : data = 16'h427A;
10'h01A8 : data = 16'h41CE;
10'h01A9 : data = 16'h4121;
10'h01AA : data = 16'h4073;
10'h01AB : data = 16'h3FC5;
10'h01AC : data = 16'h3F17;
10'h01AD : data = 16'h3E68;
10'h01AE : data = 16'h3DB8;
10'h01AF : data = 16'h3D07;
10'h01B0 : data = 16'h3C56;
10'h01B1 : data = 16'h3BA5;
10'h01B2 : data = 16'h3AF2;
10'h01B3 : data = 16'h3A40;
10'h01B4 : data = 16'h398C;
10'h01B5 : data = 16'h38D9;
10'h01B6 : data = 16'h3824;
10'h01B7 : data = 16'h376F;
10'h01B8 : data = 16'h36BA;
10'h01B9 : data = 16'h3604;
10'h01BA : data = 16'h354D;
10'h01BB : data = 16'h3496;
10'h01BC : data = 16'h33DF;
10'h01BD : data = 16'h3326;
10'h01BE : data = 16'h326E;
10'h01BF : data = 16'h31B5;
10'h01C0 : data = 16'h30FB;
10'h01C1 : data = 16'h3041;
10'h01C2 : data = 16'h2F87;
10'h01C3 : data = 16'h2ECC;
10'h01C4 : data = 16'h2E11;
10'h01C5 : data = 16'h2D55;
10'h01C6 : data = 16'h2C99;
10'h01C7 : data = 16'h2BDC;
10'h01C8 : data = 16'h2B1F;
10'h01C9 : data = 16'h2A61;
10'h01CA : data = 16'h29A3;
10'h01CB : data = 16'h28E5;
10'h01CC : data = 16'h2826;
10'h01CD : data = 16'h2767;
10'h01CE : data = 16'h26A8;
10'h01CF : data = 16'h25E8;
10'h01D0 : data = 16'h2528;
10'h01D1 : data = 16'h2467;
10'h01D2 : data = 16'h23A6;
10'h01D3 : data = 16'h22E5;
10'h01D4 : data = 16'h2223;
10'h01D5 : data = 16'h2161;
10'h01D6 : data = 16'h209F;
10'h01D7 : data = 16'h1FDD;
10'h01D8 : data = 16'h1F1A;
10'h01D9 : data = 16'h1E57;
10'h01DA : data = 16'h1D93;
10'h01DB : data = 16'h1CCF;
10'h01DC : data = 16'h1C0B;
10'h01DD : data = 16'h1B47;
10'h01DE : data = 16'h1A82;
10'h01DF : data = 16'h19BE;
10'h01E0 : data = 16'h18F9;
10'h01E1 : data = 16'h1833;
10'h01E2 : data = 16'h176E;
10'h01E3 : data = 16'h16A8;
10'h01E4 : data = 16'h15E2;
10'h01E5 : data = 16'h151C;
10'h01E6 : data = 16'h1455;
10'h01E7 : data = 16'h138F;
10'h01E8 : data = 16'h12C8;
10'h01E9 : data = 16'h1201;
10'h01EA : data = 16'h113A;
10'h01EB : data = 16'h1072;
10'h01EC : data = 16'h0FAB;
10'h01ED : data = 16'h0EE3;
10'h01EE : data = 16'h0E1C;
10'h01EF : data = 16'h0D54;
10'h01F0 : data = 16'h0C8C;
10'h01F1 : data = 16'h0BC4;
10'h01F2 : data = 16'h0AFB;
10'h01F3 : data = 16'h0A33;
10'h01F4 : data = 16'h096A;
10'h01F5 : data = 16'h08A2;
10'h01F6 : data = 16'h07D9;
10'h01F7 : data = 16'h0711;
10'h01F8 : data = 16'h0648;
10'h01F9 : data = 16'h057F;
10'h01FA : data = 16'h04B6;
10'h01FB : data = 16'h03ED;
10'h01FC : data = 16'h0324;
10'h01FD : data = 16'h025B;
10'h01FE : data = 16'h0192;
10'h01FF : data = 16'h00C9;
10'h0200 : data = 16'h0000;
10'h0201 : data = 16'hFF37;
10'h0202 : data = 16'hFE6E;
10'h0203 : data = 16'hFDA5;
10'h0204 : data = 16'hFCDC;
10'h0205 : data = 16'hFC13;
10'h0206 : data = 16'hFB4A;
10'h0207 : data = 16'hFA81;
10'h0208 : data = 16'hF9B8;
10'h0209 : data = 16'hF8EF;
10'h020A : data = 16'hF827;
10'h020B : data = 16'hF75E;
10'h020C : data = 16'hF696;
10'h020D : data = 16'hF5CD;
10'h020E : data = 16'hF505;
10'h020F : data = 16'hF43C;
10'h0210 : data = 16'hF374;
10'h0211 : data = 16'hF2AC;
10'h0212 : data = 16'hF1E4;
10'h0213 : data = 16'hF11D;
10'h0214 : data = 16'hF055;
10'h0215 : data = 16'hEF8E;
10'h0216 : data = 16'hEEC6;
10'h0217 : data = 16'hEDFF;
10'h0218 : data = 16'hED38;
10'h0219 : data = 16'hEC71;
10'h021A : data = 16'hEBAB;
10'h021B : data = 16'hEAE4;
10'h021C : data = 16'hEA1E;
10'h021D : data = 16'hE958;
10'h021E : data = 16'hE892;
10'h021F : data = 16'hE7CD;
10'h0220 : data = 16'hE707;
10'h0221 : data = 16'hE642;
10'h0222 : data = 16'hE57E;
10'h0223 : data = 16'hE4B9;
10'h0224 : data = 16'hE3F5;
10'h0225 : data = 16'hE331;
10'h0226 : data = 16'hE26D;
10'h0227 : data = 16'hE1A9;
10'h0228 : data = 16'hE0E6;
10'h0229 : data = 16'hE023;
10'h022A : data = 16'hDF61;
10'h022B : data = 16'hDE9F;
10'h022C : data = 16'hDDDD;
10'h022D : data = 16'hDD1B;
10'h022E : data = 16'hDC5A;
10'h022F : data = 16'hDB99;
10'h0230 : data = 16'hDAD8;
10'h0231 : data = 16'hDA18;
10'h0232 : data = 16'hD958;
10'h0233 : data = 16'hD899;
10'h0234 : data = 16'hD7DA;
10'h0235 : data = 16'hD71B;
10'h0236 : data = 16'hD65D;
10'h0237 : data = 16'hD59F;
10'h0238 : data = 16'hD4E1;
10'h0239 : data = 16'hD424;
10'h023A : data = 16'hD367;
10'h023B : data = 16'hD2AB;
10'h023C : data = 16'hD1EF;
10'h023D : data = 16'hD134;
10'h023E : data = 16'hD079;
10'h023F : data = 16'hCFBF;
10'h0240 : data = 16'hCF05;
10'h0241 : data = 16'hCE4B;
10'h0242 : data = 16'hCD92;
10'h0243 : data = 16'hCCDA;
10'h0244 : data = 16'hCC21;
10'h0245 : data = 16'hCB6A;
10'h0246 : data = 16'hCAB3;
10'h0247 : data = 16'hC9FC;
10'h0248 : data = 16'hC946;
10'h0249 : data = 16'hC891;
10'h024A : data = 16'hC7DC;
10'h024B : data = 16'hC727;
10'h024C : data = 16'hC674;
10'h024D : data = 16'hC5C0;
10'h024E : data = 16'hC50E;
10'h024F : data = 16'hC45B;
10'h0250 : data = 16'hC3AA;
10'h0251 : data = 16'hC2F9;
10'h0252 : data = 16'hC248;
10'h0253 : data = 16'hC198;
10'h0254 : data = 16'hC0E9;
10'h0255 : data = 16'hC03B;
10'h0256 : data = 16'hBF8D;
10'h0257 : data = 16'hBEDF;
10'h0258 : data = 16'hBE32;
10'h0259 : data = 16'hBD86;
10'h025A : data = 16'hBCDB;
10'h025B : data = 16'hBC30;
10'h025C : data = 16'hBB86;
10'h025D : data = 16'hBADC;
10'h025E : data = 16'hBA33;
10'h025F : data = 16'hB98B;
10'h0260 : data = 16'hB8E4;
10'h0261 : data = 16'hB83D;
10'h0262 : data = 16'hB797;
10'h0263 : data = 16'hB6F1;
10'h0264 : data = 16'hB64C;
10'h0265 : data = 16'hB5A8;
10'h0266 : data = 16'hB505;
10'h0267 : data = 16'hB463;
10'h0268 : data = 16'hB3C1;
10'h0269 : data = 16'hB320;
10'h026A : data = 16'hB27F;
10'h026B : data = 16'hB1E0;
10'h026C : data = 16'hB141;
10'h026D : data = 16'hB0A3;
10'h026E : data = 16'hB005;
10'h026F : data = 16'hAF69;
10'h0270 : data = 16'hAECD;
10'h0271 : data = 16'hAE32;
10'h0272 : data = 16'hAD98;
10'h0273 : data = 16'hACFE;
10'h0274 : data = 16'hAC65;
10'h0275 : data = 16'hABCE;
10'h0276 : data = 16'hAB37;
10'h0277 : data = 16'hAAA0;
10'h0278 : data = 16'hAA0B;
10'h0279 : data = 16'hA976;
10'h027A : data = 16'hA8E3;
10'h027B : data = 16'hA850;
10'h027C : data = 16'hA7BE;
10'h027D : data = 16'hA72D;
10'h027E : data = 16'hA69C;
10'h027F : data = 16'hA60D;
10'h0280 : data = 16'hA57E;
10'h0281 : data = 16'hA4F1;
10'h0282 : data = 16'hA464;
10'h0283 : data = 16'hA3D8;
10'h0284 : data = 16'hA34D;
10'h0285 : data = 16'hA2C2;
10'h0286 : data = 16'hA239;
10'h0287 : data = 16'hA1B1;
10'h0288 : data = 16'hA129;
10'h0289 : data = 16'hA0A3;
10'h028A : data = 16'hA01D;
10'h028B : data = 16'h9F98;
10'h028C : data = 16'h9F15;
10'h028D : data = 16'h9E92;
10'h028E : data = 16'h9E10;
10'h028F : data = 16'h9D8F;
10'h0290 : data = 16'h9D0F;
10'h0291 : data = 16'h9C90;
10'h0292 : data = 16'h9C12;
10'h0293 : data = 16'h9B94;
10'h0294 : data = 16'h9B18;
10'h0295 : data = 16'h9A9D;
10'h0296 : data = 16'h9A23;
10'h0297 : data = 16'h99AA;
10'h0298 : data = 16'h9931;
10'h0299 : data = 16'h98BA;
10'h029A : data = 16'h9844;
10'h029B : data = 16'h97CE;
10'h029C : data = 16'h975A;
10'h029D : data = 16'h96E7;
10'h029E : data = 16'h9675;
10'h029F : data = 16'h9603;
10'h02A0 : data = 16'h9593;
10'h02A1 : data = 16'h9524;
10'h02A2 : data = 16'h94B6;
10'h02A3 : data = 16'h9449;
10'h02A4 : data = 16'h93DD;
10'h02A5 : data = 16'h9372;
10'h02A6 : data = 16'h9308;
10'h02A7 : data = 16'h929F;
10'h02A8 : data = 16'h9237;
10'h02A9 : data = 16'h91D0;
10'h02AA : data = 16'h916A;
10'h02AB : data = 16'h9105;
10'h02AC : data = 16'h90A2;
10'h02AD : data = 16'h903F;
10'h02AE : data = 16'h8FDE;
10'h02AF : data = 16'h8F7D;
10'h02B0 : data = 16'h8F1E;
10'h02B1 : data = 16'h8EC0;
10'h02B2 : data = 16'h8E63;
10'h02B3 : data = 16'h8E07;
10'h02B4 : data = 16'h8DAC;
10'h02B5 : data = 16'h8D52;
10'h02B6 : data = 16'h8CF9;
10'h02B7 : data = 16'h8CA2;
10'h02B8 : data = 16'h8C4B;
10'h02B9 : data = 16'h8BF6;
10'h02BA : data = 16'h8BA1;
10'h02BB : data = 16'h8B4E;
10'h02BC : data = 16'h8AFC;
10'h02BD : data = 16'h8AAB;
10'h02BE : data = 16'h8A5B;
10'h02BF : data = 16'h8A0D;
10'h02C0 : data = 16'h89BF;
10'h02C1 : data = 16'h8973;
10'h02C2 : data = 16'h8928;
10'h02C3 : data = 16'h88DE;
10'h02C4 : data = 16'h8895;
10'h02C5 : data = 16'h884D;
10'h02C6 : data = 16'h8806;
10'h02C7 : data = 16'h87C1;
10'h02C8 : data = 16'h877C;
10'h02C9 : data = 16'h8739;
10'h02CA : data = 16'h86F7;
10'h02CB : data = 16'h86B6;
10'h02CC : data = 16'h8677;
10'h02CD : data = 16'h8638;
10'h02CE : data = 16'h85FB;
10'h02CF : data = 16'h85BF;
10'h02D0 : data = 16'h8584;
10'h02D1 : data = 16'h854A;
10'h02D2 : data = 16'h8512;
10'h02D3 : data = 16'h84DA;
10'h02D4 : data = 16'h84A4;
10'h02D5 : data = 16'h846F;
10'h02D6 : data = 16'h843B;
10'h02D7 : data = 16'h8408;
10'h02D8 : data = 16'h83D7;
10'h02D9 : data = 16'h83A7;
10'h02DA : data = 16'h8378;
10'h02DB : data = 16'h834A;
10'h02DC : data = 16'h831D;
10'h02DD : data = 16'h82F2;
10'h02DE : data = 16'h82C7;
10'h02DF : data = 16'h829E;
10'h02E0 : data = 16'h8277;
10'h02E1 : data = 16'h8250;
10'h02E2 : data = 16'h822B;
10'h02E3 : data = 16'h8206;
10'h02E4 : data = 16'h81E3;
10'h02E5 : data = 16'h81C2;
10'h02E6 : data = 16'h81A1;
10'h02E7 : data = 16'h8182;
10'h02E8 : data = 16'h8164;
10'h02E9 : data = 16'h8147;
10'h02EA : data = 16'h812B;
10'h02EB : data = 16'h8111;
10'h02EC : data = 16'h80F7;
10'h02ED : data = 16'h80DF;
10'h02EE : data = 16'h80C9;
10'h02EF : data = 16'h80B3;
10'h02F0 : data = 16'h809F;
10'h02F1 : data = 16'h808C;
10'h02F2 : data = 16'h807A;
10'h02F3 : data = 16'h8069;
10'h02F4 : data = 16'h805A;
10'h02F5 : data = 16'h804C;
10'h02F6 : data = 16'h803F;
10'h02F7 : data = 16'h8033;
10'h02F8 : data = 16'h8028;
10'h02F9 : data = 16'h801F;
10'h02FA : data = 16'h8017;
10'h02FB : data = 16'h8010;
10'h02FC : data = 16'h800B;
10'h02FD : data = 16'h8007;
10'h02FE : data = 16'h8003;
10'h02FF : data = 16'h8002;
10'h0300 : data = 16'h8001;
10'h0301 : data = 16'h8002;
10'h0302 : data = 16'h8003;
10'h0303 : data = 16'h8007;
10'h0304 : data = 16'h800B;
10'h0305 : data = 16'h8010;
10'h0306 : data = 16'h8017;
10'h0307 : data = 16'h801F;
10'h0308 : data = 16'h8028;
10'h0309 : data = 16'h8033;
10'h030A : data = 16'h803F;
10'h030B : data = 16'h804C;
10'h030C : data = 16'h805A;
10'h030D : data = 16'h8069;
10'h030E : data = 16'h807A;
10'h030F : data = 16'h808C;
10'h0310 : data = 16'h809F;
10'h0311 : data = 16'h80B3;
10'h0312 : data = 16'h80C9;
10'h0313 : data = 16'h80DF;
10'h0314 : data = 16'h80F7;
10'h0315 : data = 16'h8111;
10'h0316 : data = 16'h812B;
10'h0317 : data = 16'h8147;
10'h0318 : data = 16'h8164;
10'h0319 : data = 16'h8182;
10'h031A : data = 16'h81A1;
10'h031B : data = 16'h81C2;
10'h031C : data = 16'h81E3;
10'h031D : data = 16'h8206;
10'h031E : data = 16'h822B;
10'h031F : data = 16'h8250;
10'h0320 : data = 16'h8277;
10'h0321 : data = 16'h829E;
10'h0322 : data = 16'h82C7;
10'h0323 : data = 16'h82F2;
10'h0324 : data = 16'h831D;
10'h0325 : data = 16'h834A;
10'h0326 : data = 16'h8378;
10'h0327 : data = 16'h83A7;
10'h0328 : data = 16'h83D7;
10'h0329 : data = 16'h8408;
10'h032A : data = 16'h843B;
10'h032B : data = 16'h846F;
10'h032C : data = 16'h84A4;
10'h032D : data = 16'h84DA;
10'h032E : data = 16'h8512;
10'h032F : data = 16'h854A;
10'h0330 : data = 16'h8584;
10'h0331 : data = 16'h85BF;
10'h0332 : data = 16'h85FB;
10'h0333 : data = 16'h8638;
10'h0334 : data = 16'h8677;
10'h0335 : data = 16'h86B6;
10'h0336 : data = 16'h86F7;
10'h0337 : data = 16'h8739;
10'h0338 : data = 16'h877C;
10'h0339 : data = 16'h87C1;
10'h033A : data = 16'h8806;
10'h033B : data = 16'h884D;
10'h033C : data = 16'h8895;
10'h033D : data = 16'h88DE;
10'h033E : data = 16'h8928;
10'h033F : data = 16'h8973;
10'h0340 : data = 16'h89BF;
10'h0341 : data = 16'h8A0D;
10'h0342 : data = 16'h8A5B;
10'h0343 : data = 16'h8AAB;
10'h0344 : data = 16'h8AFC;
10'h0345 : data = 16'h8B4E;
10'h0346 : data = 16'h8BA1;
10'h0347 : data = 16'h8BF6;
10'h0348 : data = 16'h8C4B;
10'h0349 : data = 16'h8CA2;
10'h034A : data = 16'h8CF9;
10'h034B : data = 16'h8D52;
10'h034C : data = 16'h8DAC;
10'h034D : data = 16'h8E07;
10'h034E : data = 16'h8E63;
10'h034F : data = 16'h8EC0;
10'h0350 : data = 16'h8F1E;
10'h0351 : data = 16'h8F7D;
10'h0352 : data = 16'h8FDE;
10'h0353 : data = 16'h903F;
10'h0354 : data = 16'h90A2;
10'h0355 : data = 16'h9105;
10'h0356 : data = 16'h916A;
10'h0357 : data = 16'h91D0;
10'h0358 : data = 16'h9237;
10'h0359 : data = 16'h929F;
10'h035A : data = 16'h9308;
10'h035B : data = 16'h9372;
10'h035C : data = 16'h93DD;
10'h035D : data = 16'h9449;
10'h035E : data = 16'h94B6;
10'h035F : data = 16'h9524;
10'h0360 : data = 16'h9593;
10'h0361 : data = 16'h9603;
10'h0362 : data = 16'h9675;
10'h0363 : data = 16'h96E7;
10'h0364 : data = 16'h975A;
10'h0365 : data = 16'h97CE;
10'h0366 : data = 16'h9844;
10'h0367 : data = 16'h98BA;
10'h0368 : data = 16'h9931;
10'h0369 : data = 16'h99AA;
10'h036A : data = 16'h9A23;
10'h036B : data = 16'h9A9D;
10'h036C : data = 16'h9B18;
10'h036D : data = 16'h9B94;
10'h036E : data = 16'h9C12;
10'h036F : data = 16'h9C90;
10'h0370 : data = 16'h9D0F;
10'h0371 : data = 16'h9D8F;
10'h0372 : data = 16'h9E10;
10'h0373 : data = 16'h9E92;
10'h0374 : data = 16'h9F15;
10'h0375 : data = 16'h9F98;
10'h0376 : data = 16'hA01D;
10'h0377 : data = 16'hA0A3;
10'h0378 : data = 16'hA129;
10'h0379 : data = 16'hA1B1;
10'h037A : data = 16'hA239;
10'h037B : data = 16'hA2C2;
10'h037C : data = 16'hA34D;
10'h037D : data = 16'hA3D8;
10'h037E : data = 16'hA464;
10'h037F : data = 16'hA4F1;
10'h0380 : data = 16'hA57E;
10'h0381 : data = 16'hA60D;
10'h0382 : data = 16'hA69C;
10'h0383 : data = 16'hA72D;
10'h0384 : data = 16'hA7BE;
10'h0385 : data = 16'hA850;
10'h0386 : data = 16'hA8E3;
10'h0387 : data = 16'hA976;
10'h0388 : data = 16'hAA0B;
10'h0389 : data = 16'hAAA0;
10'h038A : data = 16'hAB37;
10'h038B : data = 16'hABCE;
10'h038C : data = 16'hAC65;
10'h038D : data = 16'hACFE;
10'h038E : data = 16'hAD98;
10'h038F : data = 16'hAE32;
10'h0390 : data = 16'hAECD;
10'h0391 : data = 16'hAF69;
10'h0392 : data = 16'hB005;
10'h0393 : data = 16'hB0A3;
10'h0394 : data = 16'hB141;
10'h0395 : data = 16'hB1E0;
10'h0396 : data = 16'hB27F;
10'h0397 : data = 16'hB320;
10'h0398 : data = 16'hB3C1;
10'h0399 : data = 16'hB463;
10'h039A : data = 16'hB505;
10'h039B : data = 16'hB5A8;
10'h039C : data = 16'hB64C;
10'h039D : data = 16'hB6F1;
10'h039E : data = 16'hB797;
10'h039F : data = 16'hB83D;
10'h03A0 : data = 16'hB8E4;
10'h03A1 : data = 16'hB98B;
10'h03A2 : data = 16'hBA33;
10'h03A3 : data = 16'hBADC;
10'h03A4 : data = 16'hBB86;
10'h03A5 : data = 16'hBC30;
10'h03A6 : data = 16'hBCDB;
10'h03A7 : data = 16'hBD86;
10'h03A8 : data = 16'hBE32;
10'h03A9 : data = 16'hBEDF;
10'h03AA : data = 16'hBF8D;
10'h03AB : data = 16'hC03B;
10'h03AC : data = 16'hC0E9;
10'h03AD : data = 16'hC198;
10'h03AE : data = 16'hC248;
10'h03AF : data = 16'hC2F9;
10'h03B0 : data = 16'hC3AA;
10'h03B1 : data = 16'hC45B;
10'h03B2 : data = 16'hC50E;
10'h03B3 : data = 16'hC5C0;
10'h03B4 : data = 16'hC674;
10'h03B5 : data = 16'hC727;
10'h03B6 : data = 16'hC7DC;
10'h03B7 : data = 16'hC891;
10'h03B8 : data = 16'hC946;
10'h03B9 : data = 16'hC9FC;
10'h03BA : data = 16'hCAB3;
10'h03BB : data = 16'hCB6A;
10'h03BC : data = 16'hCC21;
10'h03BD : data = 16'hCCDA;
10'h03BE : data = 16'hCD92;
10'h03BF : data = 16'hCE4B;
10'h03C0 : data = 16'hCF05;
10'h03C1 : data = 16'hCFBF;
10'h03C2 : data = 16'hD079;
10'h03C3 : data = 16'hD134;
10'h03C4 : data = 16'hD1EF;
10'h03C5 : data = 16'hD2AB;
10'h03C6 : data = 16'hD367;
10'h03C7 : data = 16'hD424;
10'h03C8 : data = 16'hD4E1;
10'h03C9 : data = 16'hD59F;
10'h03CA : data = 16'hD65D;
10'h03CB : data = 16'hD71B;
10'h03CC : data = 16'hD7DA;
10'h03CD : data = 16'hD899;
10'h03CE : data = 16'hD958;
10'h03CF : data = 16'hDA18;
10'h03D0 : data = 16'hDAD8;
10'h03D1 : data = 16'hDB99;
10'h03D2 : data = 16'hDC5A;
10'h03D3 : data = 16'hDD1B;
10'h03D4 : data = 16'hDDDD;
10'h03D5 : data = 16'hDE9F;
10'h03D6 : data = 16'hDF61;
10'h03D7 : data = 16'hE023;
10'h03D8 : data = 16'hE0E6;
10'h03D9 : data = 16'hE1A9;
10'h03DA : data = 16'hE26D;
10'h03DB : data = 16'hE331;
10'h03DC : data = 16'hE3F5;
10'h03DD : data = 16'hE4B9;
10'h03DE : data = 16'hE57E;
10'h03DF : data = 16'hE642;
10'h03E0 : data = 16'hE707;
10'h03E1 : data = 16'hE7CD;
10'h03E2 : data = 16'hE892;
10'h03E3 : data = 16'hE958;
10'h03E4 : data = 16'hEA1E;
10'h03E5 : data = 16'hEAE4;
10'h03E6 : data = 16'hEBAB;
10'h03E7 : data = 16'hEC71;
10'h03E8 : data = 16'hED38;
10'h03E9 : data = 16'hEDFF;
10'h03EA : data = 16'hEEC6;
10'h03EB : data = 16'hEF8E;
10'h03EC : data = 16'hF055;
10'h03ED : data = 16'hF11D;
10'h03EE : data = 16'hF1E4;
10'h03EF : data = 16'hF2AC;
10'h03F0 : data = 16'hF374;
10'h03F1 : data = 16'hF43C;
10'h03F2 : data = 16'hF505;
10'h03F3 : data = 16'hF5CD;
10'h03F4 : data = 16'hF696;
10'h03F5 : data = 16'hF75E;
10'h03F6 : data = 16'hF827;
10'h03F7 : data = 16'hF8EF;
10'h03F8 : data = 16'hF9B8;
10'h03F9 : data = 16'hFA81;
10'h03FA : data = 16'hFB4A;
10'h03FB : data = 16'hFC13;
10'h03FC : data = 16'hFCDC;
10'h03FD : data = 16'hFDA5;
10'h03FE : data = 16'hFE6E;
10'h03FF : data = 16'hFF37;


endcase
end
endmodule

