//Sine wave lookup table with 1024 points
//Regenerate using sine_wave_rom_gen.m

import opo_package::*;

module sine_lut(
 input wire [sine_lut_width-1:0] addr,
output reg [word_width-1:0] data
);

always @ * begin

case(addr)

10'h000 : data = 16'h0000;
10'h001 : data = 16'h00C9;
10'h002 : data = 16'h0192;
10'h003 : data = 16'h025B;
10'h004 : data = 16'h0324;
10'h005 : data = 16'h03ED;
10'h006 : data = 16'h04B6;
10'h007 : data = 16'h057F;
10'h008 : data = 16'h0648;
10'h009 : data = 16'h0711;
10'h00A : data = 16'h07D9;
10'h00B : data = 16'h08A2;
10'h00C : data = 16'h096A;
10'h00D : data = 16'h0A33;
10'h00E : data = 16'h0AFB;
10'h00F : data = 16'h0BC4;
10'h010 : data = 16'h0C8C;
10'h011 : data = 16'h0D54;
10'h012 : data = 16'h0E1C;
10'h013 : data = 16'h0EE3;
10'h014 : data = 16'h0FAB;
10'h015 : data = 16'h1072;
10'h016 : data = 16'h113A;
10'h017 : data = 16'h1201;
10'h018 : data = 16'h12C8;
10'h019 : data = 16'h138F;
10'h01A : data = 16'h1455;
10'h01B : data = 16'h151C;
10'h01C : data = 16'h15E2;
10'h01D : data = 16'h16A8;
10'h01E : data = 16'h176E;
10'h01F : data = 16'h1833;
10'h020 : data = 16'h18F9;
10'h021 : data = 16'h19BE;
10'h022 : data = 16'h1A82;
10'h023 : data = 16'h1B47;
10'h024 : data = 16'h1C0B;
10'h025 : data = 16'h1CCF;
10'h026 : data = 16'h1D93;
10'h027 : data = 16'h1E57;
10'h028 : data = 16'h1F1A;
10'h029 : data = 16'h1FDD;
10'h02A : data = 16'h209F;
10'h02B : data = 16'h2161;
10'h02C : data = 16'h2223;
10'h02D : data = 16'h22E5;
10'h02E : data = 16'h23A6;
10'h02F : data = 16'h2467;
10'h030 : data = 16'h2528;
10'h031 : data = 16'h25E8;
10'h032 : data = 16'h26A8;
10'h033 : data = 16'h2767;
10'h034 : data = 16'h2826;
10'h035 : data = 16'h28E5;
10'h036 : data = 16'h29A3;
10'h037 : data = 16'h2A61;
10'h038 : data = 16'h2B1F;
10'h039 : data = 16'h2BDC;
10'h03A : data = 16'h2C99;
10'h03B : data = 16'h2D55;
10'h03C : data = 16'h2E11;
10'h03D : data = 16'h2ECC;
10'h03E : data = 16'h2F87;
10'h03F : data = 16'h3041;
10'h040 : data = 16'h30FB;
10'h041 : data = 16'h31B5;
10'h042 : data = 16'h326E;
10'h043 : data = 16'h3326;
10'h044 : data = 16'h33DF;
10'h045 : data = 16'h3496;
10'h046 : data = 16'h354D;
10'h047 : data = 16'h3604;
10'h048 : data = 16'h36BA;
10'h049 : data = 16'h376F;
10'h04A : data = 16'h3824;
10'h04B : data = 16'h38D9;
10'h04C : data = 16'h398C;
10'h04D : data = 16'h3A40;
10'h04E : data = 16'h3AF2;
10'h04F : data = 16'h3BA5;
10'h050 : data = 16'h3C56;
10'h051 : data = 16'h3D07;
10'h052 : data = 16'h3DB8;
10'h053 : data = 16'h3E68;
10'h054 : data = 16'h3F17;
10'h055 : data = 16'h3FC5;
10'h056 : data = 16'h4073;
10'h057 : data = 16'h4121;
10'h058 : data = 16'h41CE;
10'h059 : data = 16'h427A;
10'h05A : data = 16'h4325;
10'h05B : data = 16'h43D0;
10'h05C : data = 16'h447A;
10'h05D : data = 16'h4524;
10'h05E : data = 16'h45CD;
10'h05F : data = 16'h4675;
10'h060 : data = 16'h471C;
10'h061 : data = 16'h47C3;
10'h062 : data = 16'h4869;
10'h063 : data = 16'h490F;
10'h064 : data = 16'h49B4;
10'h065 : data = 16'h4A58;
10'h066 : data = 16'h4AFB;
10'h067 : data = 16'h4B9D;
10'h068 : data = 16'h4C3F;
10'h069 : data = 16'h4CE0;
10'h06A : data = 16'h4D81;
10'h06B : data = 16'h4E20;
10'h06C : data = 16'h4EBF;
10'h06D : data = 16'h4F5D;
10'h06E : data = 16'h4FFB;
10'h06F : data = 16'h5097;
10'h070 : data = 16'h5133;
10'h071 : data = 16'h51CE;
10'h072 : data = 16'h5268;
10'h073 : data = 16'h5302;
10'h074 : data = 16'h539B;
10'h075 : data = 16'h5432;
10'h076 : data = 16'h54C9;
10'h077 : data = 16'h5560;
10'h078 : data = 16'h55F5;
10'h079 : data = 16'h568A;
10'h07A : data = 16'h571D;
10'h07B : data = 16'h57B0;
10'h07C : data = 16'h5842;
10'h07D : data = 16'h58D3;
10'h07E : data = 16'h5964;
10'h07F : data = 16'h59F3;
10'h080 : data = 16'h5A82;
10'h081 : data = 16'h5B0F;
10'h082 : data = 16'h5B9C;
10'h083 : data = 16'h5C28;
10'h084 : data = 16'h5CB3;
10'h085 : data = 16'h5D3E;
10'h086 : data = 16'h5DC7;
10'h087 : data = 16'h5E4F;
10'h088 : data = 16'h5ED7;
10'h089 : data = 16'h5F5D;
10'h08A : data = 16'h5FE3;
10'h08B : data = 16'h6068;
10'h08C : data = 16'h60EB;
10'h08D : data = 16'h616E;
10'h08E : data = 16'h61F0;
10'h08F : data = 16'h6271;
10'h090 : data = 16'h62F1;
10'h091 : data = 16'h6370;
10'h092 : data = 16'h63EE;
10'h093 : data = 16'h646C;
10'h094 : data = 16'h64E8;
10'h095 : data = 16'h6563;
10'h096 : data = 16'h65DD;
10'h097 : data = 16'h6656;
10'h098 : data = 16'h66CF;
10'h099 : data = 16'h6746;
10'h09A : data = 16'h67BC;
10'h09B : data = 16'h6832;
10'h09C : data = 16'h68A6;
10'h09D : data = 16'h6919;
10'h09E : data = 16'h698B;
10'h09F : data = 16'h69FD;
10'h0A0 : data = 16'h6A6D;
10'h0A1 : data = 16'h6ADC;
10'h0A2 : data = 16'h6B4A;
10'h0A3 : data = 16'h6BB7;
10'h0A4 : data = 16'h6C23;
10'h0A5 : data = 16'h6C8E;
10'h0A6 : data = 16'h6CF8;
10'h0A7 : data = 16'h6D61;
10'h0A8 : data = 16'h6DC9;
10'h0A9 : data = 16'h6E30;
10'h0AA : data = 16'h6E96;
10'h0AB : data = 16'h6EFB;
10'h0AC : data = 16'h6F5E;
10'h0AD : data = 16'h6FC1;
10'h0AE : data = 16'h7022;
10'h0AF : data = 16'h7083;
10'h0B0 : data = 16'h70E2;
10'h0B1 : data = 16'h7140;
10'h0B2 : data = 16'h719D;
10'h0B3 : data = 16'h71F9;
10'h0B4 : data = 16'h7254;
10'h0B5 : data = 16'h72AE;
10'h0B6 : data = 16'h7307;
10'h0B7 : data = 16'h735E;
10'h0B8 : data = 16'h73B5;
10'h0B9 : data = 16'h740A;
10'h0BA : data = 16'h745F;
10'h0BB : data = 16'h74B2;
10'h0BC : data = 16'h7504;
10'h0BD : data = 16'h7555;
10'h0BE : data = 16'h75A5;
10'h0BF : data = 16'h75F3;
10'h0C0 : data = 16'h7641;
10'h0C1 : data = 16'h768D;
10'h0C2 : data = 16'h76D8;
10'h0C3 : data = 16'h7722;
10'h0C4 : data = 16'h776B;
10'h0C5 : data = 16'h77B3;
10'h0C6 : data = 16'h77FA;
10'h0C7 : data = 16'h783F;
10'h0C8 : data = 16'h7884;
10'h0C9 : data = 16'h78C7;
10'h0CA : data = 16'h7909;
10'h0CB : data = 16'h794A;
10'h0CC : data = 16'h7989;
10'h0CD : data = 16'h79C8;
10'h0CE : data = 16'h7A05;
10'h0CF : data = 16'h7A41;
10'h0D0 : data = 16'h7A7C;
10'h0D1 : data = 16'h7AB6;
10'h0D2 : data = 16'h7AEE;
10'h0D3 : data = 16'h7B26;
10'h0D4 : data = 16'h7B5C;
10'h0D5 : data = 16'h7B91;
10'h0D6 : data = 16'h7BC5;
10'h0D7 : data = 16'h7BF8;
10'h0D8 : data = 16'h7C29;
10'h0D9 : data = 16'h7C59;
10'h0DA : data = 16'h7C88;
10'h0DB : data = 16'h7CB6;
10'h0DC : data = 16'h7CE3;
10'h0DD : data = 16'h7D0E;
10'h0DE : data = 16'h7D39;
10'h0DF : data = 16'h7D62;
10'h0E0 : data = 16'h7D89;
10'h0E1 : data = 16'h7DB0;
10'h0E2 : data = 16'h7DD5;
10'h0E3 : data = 16'h7DFA;
10'h0E4 : data = 16'h7E1D;
10'h0E5 : data = 16'h7E3E;
10'h0E6 : data = 16'h7E5F;
10'h0E7 : data = 16'h7E7E;
10'h0E8 : data = 16'h7E9C;
10'h0E9 : data = 16'h7EB9;
10'h0EA : data = 16'h7ED5;
10'h0EB : data = 16'h7EEF;
10'h0EC : data = 16'h7F09;
10'h0ED : data = 16'h7F21;
10'h0EE : data = 16'h7F37;
10'h0EF : data = 16'h7F4D;
10'h0F0 : data = 16'h7F61;
10'h0F1 : data = 16'h7F74;
10'h0F2 : data = 16'h7F86;
10'h0F3 : data = 16'h7F97;
10'h0F4 : data = 16'h7FA6;
10'h0F5 : data = 16'h7FB4;
10'h0F6 : data = 16'h7FC1;
10'h0F7 : data = 16'h7FCD;
10'h0F8 : data = 16'h7FD8;
10'h0F9 : data = 16'h7FE1;
10'h0FA : data = 16'h7FE9;
10'h0FB : data = 16'h7FF0;
10'h0FC : data = 16'h7FF5;
10'h0FD : data = 16'h7FF9;
10'h0FE : data = 16'h7FFD;
10'h0FF : data = 16'h7FFE;
10'h100 : data = 16'h7FFF;
10'h101 : data = 16'h7FFE;
10'h102 : data = 16'h7FFD;
10'h103 : data = 16'h7FF9;
10'h104 : data = 16'h7FF5;
10'h105 : data = 16'h7FF0;
10'h106 : data = 16'h7FE9;
10'h107 : data = 16'h7FE1;
10'h108 : data = 16'h7FD8;
10'h109 : data = 16'h7FCD;
10'h10A : data = 16'h7FC1;
10'h10B : data = 16'h7FB4;
10'h10C : data = 16'h7FA6;
10'h10D : data = 16'h7F97;
10'h10E : data = 16'h7F86;
10'h10F : data = 16'h7F74;
10'h110 : data = 16'h7F61;
10'h111 : data = 16'h7F4D;
10'h112 : data = 16'h7F37;
10'h113 : data = 16'h7F21;
10'h114 : data = 16'h7F09;
10'h115 : data = 16'h7EEF;
10'h116 : data = 16'h7ED5;
10'h117 : data = 16'h7EB9;
10'h118 : data = 16'h7E9C;
10'h119 : data = 16'h7E7E;
10'h11A : data = 16'h7E5F;
10'h11B : data = 16'h7E3E;
10'h11C : data = 16'h7E1D;
10'h11D : data = 16'h7DFA;
10'h11E : data = 16'h7DD5;
10'h11F : data = 16'h7DB0;
10'h120 : data = 16'h7D89;
10'h121 : data = 16'h7D62;
10'h122 : data = 16'h7D39;
10'h123 : data = 16'h7D0E;
10'h124 : data = 16'h7CE3;
10'h125 : data = 16'h7CB6;
10'h126 : data = 16'h7C88;
10'h127 : data = 16'h7C59;
10'h128 : data = 16'h7C29;
10'h129 : data = 16'h7BF8;
10'h12A : data = 16'h7BC5;
10'h12B : data = 16'h7B91;
10'h12C : data = 16'h7B5C;
10'h12D : data = 16'h7B26;
10'h12E : data = 16'h7AEE;
10'h12F : data = 16'h7AB6;
10'h130 : data = 16'h7A7C;
10'h131 : data = 16'h7A41;
10'h132 : data = 16'h7A05;
10'h133 : data = 16'h79C8;
10'h134 : data = 16'h7989;
10'h135 : data = 16'h794A;
10'h136 : data = 16'h7909;
10'h137 : data = 16'h78C7;
10'h138 : data = 16'h7884;
10'h139 : data = 16'h783F;
10'h13A : data = 16'h77FA;
10'h13B : data = 16'h77B3;
10'h13C : data = 16'h776B;
10'h13D : data = 16'h7722;
10'h13E : data = 16'h76D8;
10'h13F : data = 16'h768D;
10'h140 : data = 16'h7641;
10'h141 : data = 16'h75F3;
10'h142 : data = 16'h75A5;
10'h143 : data = 16'h7555;
10'h144 : data = 16'h7504;
10'h145 : data = 16'h74B2;
10'h146 : data = 16'h745F;
10'h147 : data = 16'h740A;
10'h148 : data = 16'h73B5;
10'h149 : data = 16'h735E;
10'h14A : data = 16'h7307;
10'h14B : data = 16'h72AE;
10'h14C : data = 16'h7254;
10'h14D : data = 16'h71F9;
10'h14E : data = 16'h719D;
10'h14F : data = 16'h7140;
10'h150 : data = 16'h70E2;
10'h151 : data = 16'h7083;
10'h152 : data = 16'h7022;
10'h153 : data = 16'h6FC1;
10'h154 : data = 16'h6F5E;
10'h155 : data = 16'h6EFB;
10'h156 : data = 16'h6E96;
10'h157 : data = 16'h6E30;
10'h158 : data = 16'h6DC9;
10'h159 : data = 16'h6D61;
10'h15A : data = 16'h6CF8;
10'h15B : data = 16'h6C8E;
10'h15C : data = 16'h6C23;
10'h15D : data = 16'h6BB7;
10'h15E : data = 16'h6B4A;
10'h15F : data = 16'h6ADC;
10'h160 : data = 16'h6A6D;
10'h161 : data = 16'h69FD;
10'h162 : data = 16'h698B;
10'h163 : data = 16'h6919;
10'h164 : data = 16'h68A6;
10'h165 : data = 16'h6832;
10'h166 : data = 16'h67BC;
10'h167 : data = 16'h6746;
10'h168 : data = 16'h66CF;
10'h169 : data = 16'h6656;
10'h16A : data = 16'h65DD;
10'h16B : data = 16'h6563;
10'h16C : data = 16'h64E8;
10'h16D : data = 16'h646C;
10'h16E : data = 16'h63EE;
10'h16F : data = 16'h6370;
10'h170 : data = 16'h62F1;
10'h171 : data = 16'h6271;
10'h172 : data = 16'h61F0;
10'h173 : data = 16'h616E;
10'h174 : data = 16'h60EB;
10'h175 : data = 16'h6068;
10'h176 : data = 16'h5FE3;
10'h177 : data = 16'h5F5D;
10'h178 : data = 16'h5ED7;
10'h179 : data = 16'h5E4F;
10'h17A : data = 16'h5DC7;
10'h17B : data = 16'h5D3E;
10'h17C : data = 16'h5CB3;
10'h17D : data = 16'h5C28;
10'h17E : data = 16'h5B9C;
10'h17F : data = 16'h5B0F;
10'h180 : data = 16'h5A82;
10'h181 : data = 16'h59F3;
10'h182 : data = 16'h5964;
10'h183 : data = 16'h58D3;
10'h184 : data = 16'h5842;
10'h185 : data = 16'h57B0;
10'h186 : data = 16'h571D;
10'h187 : data = 16'h568A;
10'h188 : data = 16'h55F5;
10'h189 : data = 16'h5560;
10'h18A : data = 16'h54C9;
10'h18B : data = 16'h5432;
10'h18C : data = 16'h539B;
10'h18D : data = 16'h5302;
10'h18E : data = 16'h5268;
10'h18F : data = 16'h51CE;
10'h190 : data = 16'h5133;
10'h191 : data = 16'h5097;
10'h192 : data = 16'h4FFB;
10'h193 : data = 16'h4F5D;
10'h194 : data = 16'h4EBF;
10'h195 : data = 16'h4E20;
10'h196 : data = 16'h4D81;
10'h197 : data = 16'h4CE0;
10'h198 : data = 16'h4C3F;
10'h199 : data = 16'h4B9D;
10'h19A : data = 16'h4AFB;
10'h19B : data = 16'h4A58;
10'h19C : data = 16'h49B4;
10'h19D : data = 16'h490F;
10'h19E : data = 16'h4869;
10'h19F : data = 16'h47C3;
10'h1A0 : data = 16'h471C;
10'h1A1 : data = 16'h4675;
10'h1A2 : data = 16'h45CD;
10'h1A3 : data = 16'h4524;
10'h1A4 : data = 16'h447A;
10'h1A5 : data = 16'h43D0;
10'h1A6 : data = 16'h4325;
10'h1A7 : data = 16'h427A;
10'h1A8 : data = 16'h41CE;
10'h1A9 : data = 16'h4121;
10'h1AA : data = 16'h4073;
10'h1AB : data = 16'h3FC5;
10'h1AC : data = 16'h3F17;
10'h1AD : data = 16'h3E68;
10'h1AE : data = 16'h3DB8;
10'h1AF : data = 16'h3D07;
10'h1B0 : data = 16'h3C56;
10'h1B1 : data = 16'h3BA5;
10'h1B2 : data = 16'h3AF2;
10'h1B3 : data = 16'h3A40;
10'h1B4 : data = 16'h398C;
10'h1B5 : data = 16'h38D9;
10'h1B6 : data = 16'h3824;
10'h1B7 : data = 16'h376F;
10'h1B8 : data = 16'h36BA;
10'h1B9 : data = 16'h3604;
10'h1BA : data = 16'h354D;
10'h1BB : data = 16'h3496;
10'h1BC : data = 16'h33DF;
10'h1BD : data = 16'h3326;
10'h1BE : data = 16'h326E;
10'h1BF : data = 16'h31B5;
10'h1C0 : data = 16'h30FB;
10'h1C1 : data = 16'h3041;
10'h1C2 : data = 16'h2F87;
10'h1C3 : data = 16'h2ECC;
10'h1C4 : data = 16'h2E11;
10'h1C5 : data = 16'h2D55;
10'h1C6 : data = 16'h2C99;
10'h1C7 : data = 16'h2BDC;
10'h1C8 : data = 16'h2B1F;
10'h1C9 : data = 16'h2A61;
10'h1CA : data = 16'h29A3;
10'h1CB : data = 16'h28E5;
10'h1CC : data = 16'h2826;
10'h1CD : data = 16'h2767;
10'h1CE : data = 16'h26A8;
10'h1CF : data = 16'h25E8;
10'h1D0 : data = 16'h2528;
10'h1D1 : data = 16'h2467;
10'h1D2 : data = 16'h23A6;
10'h1D3 : data = 16'h22E5;
10'h1D4 : data = 16'h2223;
10'h1D5 : data = 16'h2161;
10'h1D6 : data = 16'h209F;
10'h1D7 : data = 16'h1FDD;
10'h1D8 : data = 16'h1F1A;
10'h1D9 : data = 16'h1E57;
10'h1DA : data = 16'h1D93;
10'h1DB : data = 16'h1CCF;
10'h1DC : data = 16'h1C0B;
10'h1DD : data = 16'h1B47;
10'h1DE : data = 16'h1A82;
10'h1DF : data = 16'h19BE;
10'h1E0 : data = 16'h18F9;
10'h1E1 : data = 16'h1833;
10'h1E2 : data = 16'h176E;
10'h1E3 : data = 16'h16A8;
10'h1E4 : data = 16'h15E2;
10'h1E5 : data = 16'h151C;
10'h1E6 : data = 16'h1455;
10'h1E7 : data = 16'h138F;
10'h1E8 : data = 16'h12C8;
10'h1E9 : data = 16'h1201;
10'h1EA : data = 16'h113A;
10'h1EB : data = 16'h1072;
10'h1EC : data = 16'h0FAB;
10'h1ED : data = 16'h0EE3;
10'h1EE : data = 16'h0E1C;
10'h1EF : data = 16'h0D54;
10'h1F0 : data = 16'h0C8C;
10'h1F1 : data = 16'h0BC4;
10'h1F2 : data = 16'h0AFB;
10'h1F3 : data = 16'h0A33;
10'h1F4 : data = 16'h096A;
10'h1F5 : data = 16'h08A2;
10'h1F6 : data = 16'h07D9;
10'h1F7 : data = 16'h0711;
10'h1F8 : data = 16'h0648;
10'h1F9 : data = 16'h057F;
10'h1FA : data = 16'h04B6;
10'h1FB : data = 16'h03ED;
10'h1FC : data = 16'h0324;
10'h1FD : data = 16'h025B;
10'h1FE : data = 16'h0192;
10'h1FF : data = 16'h00C9;
10'h200 : data = 16'h0000;
10'h201 : data = 16'hFF37;
10'h202 : data = 16'hFE6E;
10'h203 : data = 16'hFDA5;
10'h204 : data = 16'hFCDC;
10'h205 : data = 16'hFC13;
10'h206 : data = 16'hFB4A;
10'h207 : data = 16'hFA81;
10'h208 : data = 16'hF9B8;
10'h209 : data = 16'hF8EF;
10'h20A : data = 16'hF827;
10'h20B : data = 16'hF75E;
10'h20C : data = 16'hF696;
10'h20D : data = 16'hF5CD;
10'h20E : data = 16'hF505;
10'h20F : data = 16'hF43C;
10'h210 : data = 16'hF374;
10'h211 : data = 16'hF2AC;
10'h212 : data = 16'hF1E4;
10'h213 : data = 16'hF11D;
10'h214 : data = 16'hF055;
10'h215 : data = 16'hEF8E;
10'h216 : data = 16'hEEC6;
10'h217 : data = 16'hEDFF;
10'h218 : data = 16'hED38;
10'h219 : data = 16'hEC71;
10'h21A : data = 16'hEBAB;
10'h21B : data = 16'hEAE4;
10'h21C : data = 16'hEA1E;
10'h21D : data = 16'hE958;
10'h21E : data = 16'hE892;
10'h21F : data = 16'hE7CD;
10'h220 : data = 16'hE707;
10'h221 : data = 16'hE642;
10'h222 : data = 16'hE57E;
10'h223 : data = 16'hE4B9;
10'h224 : data = 16'hE3F5;
10'h225 : data = 16'hE331;
10'h226 : data = 16'hE26D;
10'h227 : data = 16'hE1A9;
10'h228 : data = 16'hE0E6;
10'h229 : data = 16'hE023;
10'h22A : data = 16'hDF61;
10'h22B : data = 16'hDE9F;
10'h22C : data = 16'hDDDD;
10'h22D : data = 16'hDD1B;
10'h22E : data = 16'hDC5A;
10'h22F : data = 16'hDB99;
10'h230 : data = 16'hDAD8;
10'h231 : data = 16'hDA18;
10'h232 : data = 16'hD958;
10'h233 : data = 16'hD899;
10'h234 : data = 16'hD7DA;
10'h235 : data = 16'hD71B;
10'h236 : data = 16'hD65D;
10'h237 : data = 16'hD59F;
10'h238 : data = 16'hD4E1;
10'h239 : data = 16'hD424;
10'h23A : data = 16'hD367;
10'h23B : data = 16'hD2AB;
10'h23C : data = 16'hD1EF;
10'h23D : data = 16'hD134;
10'h23E : data = 16'hD079;
10'h23F : data = 16'hCFBF;
10'h240 : data = 16'hCF05;
10'h241 : data = 16'hCE4B;
10'h242 : data = 16'hCD92;
10'h243 : data = 16'hCCDA;
10'h244 : data = 16'hCC21;
10'h245 : data = 16'hCB6A;
10'h246 : data = 16'hCAB3;
10'h247 : data = 16'hC9FC;
10'h248 : data = 16'hC946;
10'h249 : data = 16'hC891;
10'h24A : data = 16'hC7DC;
10'h24B : data = 16'hC727;
10'h24C : data = 16'hC674;
10'h24D : data = 16'hC5C0;
10'h24E : data = 16'hC50E;
10'h24F : data = 16'hC45B;
10'h250 : data = 16'hC3AA;
10'h251 : data = 16'hC2F9;
10'h252 : data = 16'hC248;
10'h253 : data = 16'hC198;
10'h254 : data = 16'hC0E9;
10'h255 : data = 16'hC03B;
10'h256 : data = 16'hBF8D;
10'h257 : data = 16'hBEDF;
10'h258 : data = 16'hBE32;
10'h259 : data = 16'hBD86;
10'h25A : data = 16'hBCDB;
10'h25B : data = 16'hBC30;
10'h25C : data = 16'hBB86;
10'h25D : data = 16'hBADC;
10'h25E : data = 16'hBA33;
10'h25F : data = 16'hB98B;
10'h260 : data = 16'hB8E4;
10'h261 : data = 16'hB83D;
10'h262 : data = 16'hB797;
10'h263 : data = 16'hB6F1;
10'h264 : data = 16'hB64C;
10'h265 : data = 16'hB5A8;
10'h266 : data = 16'hB505;
10'h267 : data = 16'hB463;
10'h268 : data = 16'hB3C1;
10'h269 : data = 16'hB320;
10'h26A : data = 16'hB27F;
10'h26B : data = 16'hB1E0;
10'h26C : data = 16'hB141;
10'h26D : data = 16'hB0A3;
10'h26E : data = 16'hB005;
10'h26F : data = 16'hAF69;
10'h270 : data = 16'hAECD;
10'h271 : data = 16'hAE32;
10'h272 : data = 16'hAD98;
10'h273 : data = 16'hACFE;
10'h274 : data = 16'hAC65;
10'h275 : data = 16'hABCE;
10'h276 : data = 16'hAB37;
10'h277 : data = 16'hAAA0;
10'h278 : data = 16'hAA0B;
10'h279 : data = 16'hA976;
10'h27A : data = 16'hA8E3;
10'h27B : data = 16'hA850;
10'h27C : data = 16'hA7BE;
10'h27D : data = 16'hA72D;
10'h27E : data = 16'hA69C;
10'h27F : data = 16'hA60D;
10'h280 : data = 16'hA57E;
10'h281 : data = 16'hA4F1;
10'h282 : data = 16'hA464;
10'h283 : data = 16'hA3D8;
10'h284 : data = 16'hA34D;
10'h285 : data = 16'hA2C2;
10'h286 : data = 16'hA239;
10'h287 : data = 16'hA1B1;
10'h288 : data = 16'hA129;
10'h289 : data = 16'hA0A3;
10'h28A : data = 16'hA01D;
10'h28B : data = 16'h9F98;
10'h28C : data = 16'h9F15;
10'h28D : data = 16'h9E92;
10'h28E : data = 16'h9E10;
10'h28F : data = 16'h9D8F;
10'h290 : data = 16'h9D0F;
10'h291 : data = 16'h9C90;
10'h292 : data = 16'h9C12;
10'h293 : data = 16'h9B94;
10'h294 : data = 16'h9B18;
10'h295 : data = 16'h9A9D;
10'h296 : data = 16'h9A23;
10'h297 : data = 16'h99AA;
10'h298 : data = 16'h9931;
10'h299 : data = 16'h98BA;
10'h29A : data = 16'h9844;
10'h29B : data = 16'h97CE;
10'h29C : data = 16'h975A;
10'h29D : data = 16'h96E7;
10'h29E : data = 16'h9675;
10'h29F : data = 16'h9603;
10'h2A0 : data = 16'h9593;
10'h2A1 : data = 16'h9524;
10'h2A2 : data = 16'h94B6;
10'h2A3 : data = 16'h9449;
10'h2A4 : data = 16'h93DD;
10'h2A5 : data = 16'h9372;
10'h2A6 : data = 16'h9308;
10'h2A7 : data = 16'h929F;
10'h2A8 : data = 16'h9237;
10'h2A9 : data = 16'h91D0;
10'h2AA : data = 16'h916A;
10'h2AB : data = 16'h9105;
10'h2AC : data = 16'h90A2;
10'h2AD : data = 16'h903F;
10'h2AE : data = 16'h8FDE;
10'h2AF : data = 16'h8F7D;
10'h2B0 : data = 16'h8F1E;
10'h2B1 : data = 16'h8EC0;
10'h2B2 : data = 16'h8E63;
10'h2B3 : data = 16'h8E07;
10'h2B4 : data = 16'h8DAC;
10'h2B5 : data = 16'h8D52;
10'h2B6 : data = 16'h8CF9;
10'h2B7 : data = 16'h8CA2;
10'h2B8 : data = 16'h8C4B;
10'h2B9 : data = 16'h8BF6;
10'h2BA : data = 16'h8BA1;
10'h2BB : data = 16'h8B4E;
10'h2BC : data = 16'h8AFC;
10'h2BD : data = 16'h8AAB;
10'h2BE : data = 16'h8A5B;
10'h2BF : data = 16'h8A0D;
10'h2C0 : data = 16'h89BF;
10'h2C1 : data = 16'h8973;
10'h2C2 : data = 16'h8928;
10'h2C3 : data = 16'h88DE;
10'h2C4 : data = 16'h8895;
10'h2C5 : data = 16'h884D;
10'h2C6 : data = 16'h8806;
10'h2C7 : data = 16'h87C1;
10'h2C8 : data = 16'h877C;
10'h2C9 : data = 16'h8739;
10'h2CA : data = 16'h86F7;
10'h2CB : data = 16'h86B6;
10'h2CC : data = 16'h8677;
10'h2CD : data = 16'h8638;
10'h2CE : data = 16'h85FB;
10'h2CF : data = 16'h85BF;
10'h2D0 : data = 16'h8584;
10'h2D1 : data = 16'h854A;
10'h2D2 : data = 16'h8512;
10'h2D3 : data = 16'h84DA;
10'h2D4 : data = 16'h84A4;
10'h2D5 : data = 16'h846F;
10'h2D6 : data = 16'h843B;
10'h2D7 : data = 16'h8408;
10'h2D8 : data = 16'h83D7;
10'h2D9 : data = 16'h83A7;
10'h2DA : data = 16'h8378;
10'h2DB : data = 16'h834A;
10'h2DC : data = 16'h831D;
10'h2DD : data = 16'h82F2;
10'h2DE : data = 16'h82C7;
10'h2DF : data = 16'h829E;
10'h2E0 : data = 16'h8277;
10'h2E1 : data = 16'h8250;
10'h2E2 : data = 16'h822B;
10'h2E3 : data = 16'h8206;
10'h2E4 : data = 16'h81E3;
10'h2E5 : data = 16'h81C2;
10'h2E6 : data = 16'h81A1;
10'h2E7 : data = 16'h8182;
10'h2E8 : data = 16'h8164;
10'h2E9 : data = 16'h8147;
10'h2EA : data = 16'h812B;
10'h2EB : data = 16'h8111;
10'h2EC : data = 16'h80F7;
10'h2ED : data = 16'h80DF;
10'h2EE : data = 16'h80C9;
10'h2EF : data = 16'h80B3;
10'h2F0 : data = 16'h809F;
10'h2F1 : data = 16'h808C;
10'h2F2 : data = 16'h807A;
10'h2F3 : data = 16'h8069;
10'h2F4 : data = 16'h805A;
10'h2F5 : data = 16'h804C;
10'h2F6 : data = 16'h803F;
10'h2F7 : data = 16'h8033;
10'h2F8 : data = 16'h8028;
10'h2F9 : data = 16'h801F;
10'h2FA : data = 16'h8017;
10'h2FB : data = 16'h8010;
10'h2FC : data = 16'h800B;
10'h2FD : data = 16'h8007;
10'h2FE : data = 16'h8003;
10'h2FF : data = 16'h8002;
10'h300 : data = 16'h8001;
10'h301 : data = 16'h8002;
10'h302 : data = 16'h8003;
10'h303 : data = 16'h8007;
10'h304 : data = 16'h800B;
10'h305 : data = 16'h8010;
10'h306 : data = 16'h8017;
10'h307 : data = 16'h801F;
10'h308 : data = 16'h8028;
10'h309 : data = 16'h8033;
10'h30A : data = 16'h803F;
10'h30B : data = 16'h804C;
10'h30C : data = 16'h805A;
10'h30D : data = 16'h8069;
10'h30E : data = 16'h807A;
10'h30F : data = 16'h808C;
10'h310 : data = 16'h809F;
10'h311 : data = 16'h80B3;
10'h312 : data = 16'h80C9;
10'h313 : data = 16'h80DF;
10'h314 : data = 16'h80F7;
10'h315 : data = 16'h8111;
10'h316 : data = 16'h812B;
10'h317 : data = 16'h8147;
10'h318 : data = 16'h8164;
10'h319 : data = 16'h8182;
10'h31A : data = 16'h81A1;
10'h31B : data = 16'h81C2;
10'h31C : data = 16'h81E3;
10'h31D : data = 16'h8206;
10'h31E : data = 16'h822B;
10'h31F : data = 16'h8250;
10'h320 : data = 16'h8277;
10'h321 : data = 16'h829E;
10'h322 : data = 16'h82C7;
10'h323 : data = 16'h82F2;
10'h324 : data = 16'h831D;
10'h325 : data = 16'h834A;
10'h326 : data = 16'h8378;
10'h327 : data = 16'h83A7;
10'h328 : data = 16'h83D7;
10'h329 : data = 16'h8408;
10'h32A : data = 16'h843B;
10'h32B : data = 16'h846F;
10'h32C : data = 16'h84A4;
10'h32D : data = 16'h84DA;
10'h32E : data = 16'h8512;
10'h32F : data = 16'h854A;
10'h330 : data = 16'h8584;
10'h331 : data = 16'h85BF;
10'h332 : data = 16'h85FB;
10'h333 : data = 16'h8638;
10'h334 : data = 16'h8677;
10'h335 : data = 16'h86B6;
10'h336 : data = 16'h86F7;
10'h337 : data = 16'h8739;
10'h338 : data = 16'h877C;
10'h339 : data = 16'h87C1;
10'h33A : data = 16'h8806;
10'h33B : data = 16'h884D;
10'h33C : data = 16'h8895;
10'h33D : data = 16'h88DE;
10'h33E : data = 16'h8928;
10'h33F : data = 16'h8973;
10'h340 : data = 16'h89BF;
10'h341 : data = 16'h8A0D;
10'h342 : data = 16'h8A5B;
10'h343 : data = 16'h8AAB;
10'h344 : data = 16'h8AFC;
10'h345 : data = 16'h8B4E;
10'h346 : data = 16'h8BA1;
10'h347 : data = 16'h8BF6;
10'h348 : data = 16'h8C4B;
10'h349 : data = 16'h8CA2;
10'h34A : data = 16'h8CF9;
10'h34B : data = 16'h8D52;
10'h34C : data = 16'h8DAC;
10'h34D : data = 16'h8E07;
10'h34E : data = 16'h8E63;
10'h34F : data = 16'h8EC0;
10'h350 : data = 16'h8F1E;
10'h351 : data = 16'h8F7D;
10'h352 : data = 16'h8FDE;
10'h353 : data = 16'h903F;
10'h354 : data = 16'h90A2;
10'h355 : data = 16'h9105;
10'h356 : data = 16'h916A;
10'h357 : data = 16'h91D0;
10'h358 : data = 16'h9237;
10'h359 : data = 16'h929F;
10'h35A : data = 16'h9308;
10'h35B : data = 16'h9372;
10'h35C : data = 16'h93DD;
10'h35D : data = 16'h9449;
10'h35E : data = 16'h94B6;
10'h35F : data = 16'h9524;
10'h360 : data = 16'h9593;
10'h361 : data = 16'h9603;
10'h362 : data = 16'h9675;
10'h363 : data = 16'h96E7;
10'h364 : data = 16'h975A;
10'h365 : data = 16'h97CE;
10'h366 : data = 16'h9844;
10'h367 : data = 16'h98BA;
10'h368 : data = 16'h9931;
10'h369 : data = 16'h99AA;
10'h36A : data = 16'h9A23;
10'h36B : data = 16'h9A9D;
10'h36C : data = 16'h9B18;
10'h36D : data = 16'h9B94;
10'h36E : data = 16'h9C12;
10'h36F : data = 16'h9C90;
10'h370 : data = 16'h9D0F;
10'h371 : data = 16'h9D8F;
10'h372 : data = 16'h9E10;
10'h373 : data = 16'h9E92;
10'h374 : data = 16'h9F15;
10'h375 : data = 16'h9F98;
10'h376 : data = 16'hA01D;
10'h377 : data = 16'hA0A3;
10'h378 : data = 16'hA129;
10'h379 : data = 16'hA1B1;
10'h37A : data = 16'hA239;
10'h37B : data = 16'hA2C2;
10'h37C : data = 16'hA34D;
10'h37D : data = 16'hA3D8;
10'h37E : data = 16'hA464;
10'h37F : data = 16'hA4F1;
10'h380 : data = 16'hA57E;
10'h381 : data = 16'hA60D;
10'h382 : data = 16'hA69C;
10'h383 : data = 16'hA72D;
10'h384 : data = 16'hA7BE;
10'h385 : data = 16'hA850;
10'h386 : data = 16'hA8E3;
10'h387 : data = 16'hA976;
10'h388 : data = 16'hAA0B;
10'h389 : data = 16'hAAA0;
10'h38A : data = 16'hAB37;
10'h38B : data = 16'hABCE;
10'h38C : data = 16'hAC65;
10'h38D : data = 16'hACFE;
10'h38E : data = 16'hAD98;
10'h38F : data = 16'hAE32;
10'h390 : data = 16'hAECD;
10'h391 : data = 16'hAF69;
10'h392 : data = 16'hB005;
10'h393 : data = 16'hB0A3;
10'h394 : data = 16'hB141;
10'h395 : data = 16'hB1E0;
10'h396 : data = 16'hB27F;
10'h397 : data = 16'hB320;
10'h398 : data = 16'hB3C1;
10'h399 : data = 16'hB463;
10'h39A : data = 16'hB505;
10'h39B : data = 16'hB5A8;
10'h39C : data = 16'hB64C;
10'h39D : data = 16'hB6F1;
10'h39E : data = 16'hB797;
10'h39F : data = 16'hB83D;
10'h3A0 : data = 16'hB8E4;
10'h3A1 : data = 16'hB98B;
10'h3A2 : data = 16'hBA33;
10'h3A3 : data = 16'hBADC;
10'h3A4 : data = 16'hBB86;
10'h3A5 : data = 16'hBC30;
10'h3A6 : data = 16'hBCDB;
10'h3A7 : data = 16'hBD86;
10'h3A8 : data = 16'hBE32;
10'h3A9 : data = 16'hBEDF;
10'h3AA : data = 16'hBF8D;
10'h3AB : data = 16'hC03B;
10'h3AC : data = 16'hC0E9;
10'h3AD : data = 16'hC198;
10'h3AE : data = 16'hC248;
10'h3AF : data = 16'hC2F9;
10'h3B0 : data = 16'hC3AA;
10'h3B1 : data = 16'hC45B;
10'h3B2 : data = 16'hC50E;
10'h3B3 : data = 16'hC5C0;
10'h3B4 : data = 16'hC674;
10'h3B5 : data = 16'hC727;
10'h3B6 : data = 16'hC7DC;
10'h3B7 : data = 16'hC891;
10'h3B8 : data = 16'hC946;
10'h3B9 : data = 16'hC9FC;
10'h3BA : data = 16'hCAB3;
10'h3BB : data = 16'hCB6A;
10'h3BC : data = 16'hCC21;
10'h3BD : data = 16'hCCDA;
10'h3BE : data = 16'hCD92;
10'h3BF : data = 16'hCE4B;
10'h3C0 : data = 16'hCF05;
10'h3C1 : data = 16'hCFBF;
10'h3C2 : data = 16'hD079;
10'h3C3 : data = 16'hD134;
10'h3C4 : data = 16'hD1EF;
10'h3C5 : data = 16'hD2AB;
10'h3C6 : data = 16'hD367;
10'h3C7 : data = 16'hD424;
10'h3C8 : data = 16'hD4E1;
10'h3C9 : data = 16'hD59F;
10'h3CA : data = 16'hD65D;
10'h3CB : data = 16'hD71B;
10'h3CC : data = 16'hD7DA;
10'h3CD : data = 16'hD899;
10'h3CE : data = 16'hD958;
10'h3CF : data = 16'hDA18;
10'h3D0 : data = 16'hDAD8;
10'h3D1 : data = 16'hDB99;
10'h3D2 : data = 16'hDC5A;
10'h3D3 : data = 16'hDD1B;
10'h3D4 : data = 16'hDDDD;
10'h3D5 : data = 16'hDE9F;
10'h3D6 : data = 16'hDF61;
10'h3D7 : data = 16'hE023;
10'h3D8 : data = 16'hE0E6;
10'h3D9 : data = 16'hE1A9;
10'h3DA : data = 16'hE26D;
10'h3DB : data = 16'hE331;
10'h3DC : data = 16'hE3F5;
10'h3DD : data = 16'hE4B9;
10'h3DE : data = 16'hE57E;
10'h3DF : data = 16'hE642;
10'h3E0 : data = 16'hE707;
10'h3E1 : data = 16'hE7CD;
10'h3E2 : data = 16'hE892;
10'h3E3 : data = 16'hE958;
10'h3E4 : data = 16'hEA1E;
10'h3E5 : data = 16'hEAE4;
10'h3E6 : data = 16'hEBAB;
10'h3E7 : data = 16'hEC71;
10'h3E8 : data = 16'hED38;
10'h3E9 : data = 16'hEDFF;
10'h3EA : data = 16'hEEC6;
10'h3EB : data = 16'hEF8E;
10'h3EC : data = 16'hF055;
10'h3ED : data = 16'hF11D;
10'h3EE : data = 16'hF1E4;
10'h3EF : data = 16'hF2AC;
10'h3F0 : data = 16'hF374;
10'h3F1 : data = 16'hF43C;
10'h3F2 : data = 16'hF505;
10'h3F3 : data = 16'hF5CD;
10'h3F4 : data = 16'hF696;
10'h3F5 : data = 16'hF75E;
10'h3F6 : data = 16'hF827;
10'h3F7 : data = 16'hF8EF;
10'h3F8 : data = 16'hF9B8;
10'h3F9 : data = 16'hFA81;
10'h3FA : data = 16'hFB4A;
10'h3FB : data = 16'hFC13;
10'h3FC : data = 16'hFCDC;
10'h3FD : data = 16'hFDA5;
10'h3FE : data = 16'hFE6E;
10'h3FF : data = 16'hFF37;


endcase
end
endmodule

