package opo_package;


parameter word_width = 16;
parameter sine_lut_width = 10;
parameter config_reg_width = 128;

endpackage